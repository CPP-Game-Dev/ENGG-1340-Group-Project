1|Camping Boots|Max SP +10|0|0|10|0|0|0|0|0|0|0|0|0
2|Old Belt|Pickaxe Capacity +1|0|0|0|0|0|0|1|0|0|0|0|0
3|Hoarders Backpack|Ration Capacity +2|0|0|0|0|0|2|0|0|0|0|0|0
4|Charred Steak|Max SP +15|0|0|15|0|0|0|0|0|0|0|0|0
5|Rotten Egg|Ration Effectiveness +3|0|0|0|3|0|0|0|0|0|0|0|0
6|Oil Lamp|FOV +1|0|0|0|0|1|0|0|0|0|0|0|0
7|Expired Milk|Ration Effectiveness +1_Max SP +5|0|0|5|5|0|0|0|0|0|0|0|0
8|Worn Sneakers|Max SP +5_10% chance to not conume stamina when moving|0|1|5|0|0|0|0|0|0|0|0|0
9|Spinach Leaf|Max SP +10%|0|0|0|0|0|0|0|0.1|0|0|0|0
10|Ink Bottle|Leave ink marks behind as you move|0|1|0|0|0|0|0|0|0|0|0|0
11|Comically Oversized Cookie|Effectiveness of Rations +8|0|0|0|8|0|0|0|0|0|0|0|0
12|Mutated Potato|Ration Capacity -1_+1 Ration every 50 steps|0|1|0|0|0|0|0|0|0|0|0|0
13|Moldy Cheese|Effectiveness of Rations -25%_+20% chance to not consume Ration|0|1|0|0|0|0|0|0|0.25|0|0|0
14|Sleeping Bag|+10 SP at the end of a level|0|1|0|0|0|0|0|0|0|0|0|0
15|Camping Backpack|Pickaxe & Ration Capacity +1|1|0|0|0|0|1|1|0|0|0|0|0
16|Camping Flashlight|FOV +2|1|0|0|0|2|0|0|0|0|0|0|0
17|Charm Of Satiation|+5 SP when picking up anything_Max SP +20|1|1|20|0|0|0|0|0|0|0|0|0
18|Emergency Rations|+100% SP when it reaches 0 (once)|1|0|0|0|0|0|0|0|0|0|0|0
19|Roller Skates|Max Stamin +5_33% chance to not consume energy when moving|1|1|5|0|0|0|0|0|0|0|0|0
20|Lit Torch|FOV +3_Burns out after 150 steps|1|1|0|0|3|0|0|0|0|0|0|0
21|M.R.E.|Effectiveness of Rations +10_ Max SP +10%|1|0|10|0|0|0|0|0.1|0|0|0|0
22|Millitary Backpack|Ration Capacity +5_Effectiveness of Rations -10%|1|0|0|0|5|0|0|0|-0.1|0|0|0
23|Enchanted Bracelet|+15 SP at the end of a level|1|1|0|0|0|0|0|0|0|0|0|0
24|Guide to Underground Exploration (Vol 1)|Increase the amount of collectables by 2|1|1|0|0|0|0|0|0|0|0|0|0
25|Guide to Underground Exploration (Vol 2)|20% chance to +3 stamina every step|1|1|0|0|0|0|0|0|0|0|0|0
26|Bundle Of Breadsticks|Max SP +20%|1|0|0|0|0|0|0|0.2|0|0|0|0
27|Headlights|FOV +3|2|0|0|0|3|0|0|0|0|0|0|0
28|Telescope Glasses|FOV +75%, can no longer see yourself|2|1|0|0|0|0|0|0|0|0.75|0|0
29|Metal Detector|Chests will produce rarer items|2|1|0|0|0|0|0|0|0|0|0|0
30|Magic Mushroom|Effectiveness of Rations +50%, Max SP -33%|2|0|0|0|0|0|0|-0.33|0.5|0|0|0
31|Mining Helmet|+50% chance to not consume a Pickaxe when breaking walls|2|1|0|0|0|0|0|0|0|0|0|0
32|Suspicious Pills|Effectiveness of Rations +1 per 3 steps|2|1|0|0|0|0|0|0|0|0|0|0
33|Insulin Injection|Effectiveness of Rations +15, FOV -1|2|1|0|15|-1|0|0|0|0|0|0|0
34|Wheelchair|25% chance to not consume SP when moving|2|1|0|0|0|0|0|0|0|0|0|0
35|Hiking Staff|+1 Max SP per 5 steps , Max SP -20|2|1|-20|0|0|0|0|0|0|0|0|0
36|Premium Sportswear|Max SP +35%, Ration & Rickaxe Capacity +1|2|1|0|0|0|1|1|0.35|0|0|0|0
37|Hermes Boots|80% chance to not consume stamina when moving|3|1|0|0|0|0|0|0|0|0|0|0
38|Quadruple Espresso|SP Capacity +75%|3|0|0|0|0|0|0|0.75|0|0|0|0
39|Auringonsiemen|You can see everything|3|1|0|0|0|0|0|0|0|0|0|0
40|Alpha Star|Permanent +10 Max SP when completing a level|3|1|0|0|0|0|0|0|0|0|0|0
41|RedBull|Effect of Energy Drinks +150%|3|1|0|0|0|0|0|0|0|0|0|0