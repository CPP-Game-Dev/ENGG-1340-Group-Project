1|Camping Boots|Max Stamina +10|0|0|10|0|0|0|0|0|0|0|0|0
2|Old Belt|Pickaxe Capacity +1, Ration Capacity -1|0|0|0|0|0|-1|1|0|0|0|0|0
3|Hoarders Backpack|Ration Capacity +2|0|0|0|0|0|2|0|0|0|0|0|0
4|Charred Steak|Max Stamina +15|0|0|15|0|0|0|0|0|0|0|0|0
5|Rotten Egg|Ration Effectiveness +3|0|0|0|3|0|0|0|0|0|0|0|0
6|Oil Lamp|FOV +1|0|0|0|0|1|0|0|0|0|0|0|0
7|Expired Milk|Ration Effectiveness +1, Max Stamina +5|0|0|5|5|0|0|0|0|0|0|0|0
8|Worn Sneakers|Max Stamina +5, 10% chance to move for free|0|1|5|0|0|0|0|0|0|0|0|0
9|Spinach Leaf|Max Stamina +10%|0|0|0|0|0|0|0|0.1|0|0|0|0
10|Ink Bottle|Leave ink marks behind as you move|0|1|0|0|0|0|0|0|0|0|0|0
11|Comically Oversized Cookie|Increase effectiveness of Rations by 8|0|0|0|8|0|0|0|0|0|0|0|0
12|Mutated Potato|Decrease Ration Capacity by 1, generate 1 Ration for every 60 steps taken, increase Max Stamina by 5|0|1|5|0|0|0|0|0|0|0|0|0
13|Moldy Cheese|Decrease effectiveness of Rations by 25%, has 10% chance to not consume a Ration when eating|0|1|0|0|0|0|0|0|0.25|0|0|0
14|Sleeping Bag|Regenerate 10 additional Stamina at the end of a level|0|1|0|0|0|0|0|0|0|0|0|0
15|Camping Backpack|Increase Pickaxe & Ration Capacity by 1|1|0|0|0|0|1|1|0|0|0|0|0
16|Camping Flashlight|Increase FOV by 2|1|0|0|0|2|0|0|0|0|0|0|0
17|Charm Of Satiation|Regenerate 5 Stamina when picking up a Collectable, increase Max Stamina by 20|1|1|20|0|0|0|0|0|0|0|0|0
18|Emergency Rations|Fully regenerates Stamina when it reaches 0|1|0|0|0|0|0|0|0|0|0|0|0
19|Roller Skates|Max Stamin +5, has 33% chance to move for free|1|1|5|0|0|0|0|0|0|0|0|0
20|Lit Torch|Increase FOV by 3, burns out permanently after 150 steps|1|1|0|0|3|0|0|0|0|0|0|0
21|M.R.E.|Increase effectiveness of Rations by 10, increase Max Stamina 10%|1|0|10|0|0|0|0|0.1|0|0|0|0
22|Millitary Backpack|Increase Ration Capacity by 5, decrease effectiveness of Rations by 10%|1|0|0|0|5|0|0|0|-0.1|0|0|0
23|Enchanted Bracelet|Regenerates 15 addi Stamina at the end of a level|1|1|0|0|0|0|0|0|0|0|0|0
24|Guide to Underground Exploration (Vol 1)|Highlights the nearest Ration on the map|1|1|0|0|0|0|0|0|0|0|0|0
25|Guide to Underground Exploration (Vol 2)|Highlights the nearest Energy Drink on the map|1|1|0|0|0|0|0|0|0|0|0|0
26|Bundle Of Breadsticks|Increase Max Stamina by 20%|1|0|0|0|0|0|0|0.2|0|0|0|0
27|Headlights|Increase FOV by 3|2|0|0|0|3|0|0|0|0|0|0|0
28|Telescope Glasses|Increase FOV by 75%, can no longer see in a 3-tile radius|2|1|0|0|0|0|0|0|0|0.75|0|0
29|Metal Detector|Highlights the nearest Chest on the map|2|1|0|0|0|0|0|0|0|0|0|0
30|Magic Mushroom|Increase the effectiveness of Rations by 50%, decrease Max Stamina by 33%|2|0|0|0|0|0|0|-0.33|0.5|0|0|0
31|Mining Helmet|Has a 50% chance to not consume a Pickaxe when breaking walls|2|1|0|0|0|0|0|0|0|0|0|0
32|Suspicious Pills|Rations become Energy Drinks, you can no longer carry rations|2|1|0|0|0|0|0|0|0|0|-999|0
33|Insulin Injection|Increase the effectiveness of Rations by 15, decrease FOV by 1|2|1|0|15|-1|0|0|0|0|0|0|0
34|Wheelchair|Has a 25% chance to not consume Stamina when moving|2|1|0|0|0|0|0|0|0|0|0|0
35|Hiking Staff|Recovers 1 Stamina per 5 steps , increase Max Stamina by 10|2|1|10|0|0|0|0|0|0|0|0|0
36|Premium Sportswear|Increase Max Stamina by 35%, ration & pickaxe capacity by 1|2|1|0|0|0|1|1|0.35|0|0|0|0
37|Hermes Boots|Has an 80% chance to not consume stamina when moving|3|1|0|0|0|0|0|0|0|0|0|0
38|Quadruple Espresso|Increase Stamina Capacity by 75%|3|0|0|0|0|0|0|0.75|0|0|0|0
39|Auringonsiemen|You can now see everything|3|1|0|0|0|0|0|0|0|0|0|0
40|Alpha Star|Highlights the exit on the map|3|1|0|0|0|0|0|0|0|0|0|0